`timescale 1ns / 1ps

module tb_or;
    reg a, b;
    wire or_out;
         
    demux_or_gate dut(a, b, or_out);
    initial begin
            a= 1'b0; b= 1'b0;
        #10 a= 1'b0; b= 1'b1;
        #10 a= 1'b1; b= 1'b0;
        #10 a= 1'b1; b= 1'b1;
    end
    initial 
     begin
       $dumpfile("tb_or.vcd");
       $dumpvars(0,tb_or);
       $monitor("a: %b  b: %b  or: %b ",a, b, or_out);
     #40 $finish;
     end
endmodule
module SR_flipflop(
input clk, reset,S,R,
output reg Q
);

always@(posedge clk) begin 
if(reset) Q<=1'b0 ;

else begin 
case({S,R})
2'b00: Q<=Q;
2'b01: Q<=1'b0;
2'b10: Q<=1'b1 ;
default : Q<=2'bxx;
endcase
end
end
endmodule 
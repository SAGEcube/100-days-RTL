`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 11/02/2025 10:34:26 PM
// Design Name: 
// Module Name: test_bench
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


`timescale 1ns / 1ps

module test_bench;
reg clk,rst,J,K;
wire Q_sr, Q_d, Q_t;

  JK_using_SR_D_T dut(J, K, clk, rst, Q_sr, Q_d, Q_t);
initial begin 
        clk = 0;
       forever #5 clk = ~clk;
       end 
       
 initial begin
        rst=1;
        J = 0;
        K = 0;
        #10;
        rst=0;
    end
    
    always begin
        J=0;
        K=0;
        #10;
        J=0;
        K=1;
        #10;
        J=1;
        K=0;
        #10;
        J=1;
        K=1;
        #10;

    end
  initial begin
  $dumpfile("test_bench.vcd");
  $dumpvars(0,test_bench);
  $monitor("\t clk: %d  J: %d  K: %d  Q_sr: %d  Q_d: %d  Q_t:%d", clk,J,K,Q_sr, Q_d, Q_t);
  #90 $finish;
  end
endmodule

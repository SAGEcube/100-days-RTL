module decoder_2_4(
  input [1:0] i ,
  output reg [3:0] y);
  
  always@(*) begin 
    y = 0 ;
    case(i) 
      2'b00: y[0] = 1'b1 ;
      2'b00: y[1] = 1'b1 ;
      2'b00: y[2] = 1'b1 ;
      2'b00: y[3] = 1'b1 ;
    endcase
  end
endmodule 

module decoder_or(
  input a,b ,
  output or_g
);
  wire[3:0] w;
  decoder_2_4  orgate({a,b},w);
  
  assign or_g = ~w[0] ;
endmodule 
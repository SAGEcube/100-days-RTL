`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 11/01/2025 10:35:57 AM
// Design Name: 
// Module Name: test_bench
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////



`timescale 1ns / 1ps

module test_bench;
reg S, R, clk, rst;
wire Q_jk, Q_d, Q_t;

  SR_using_JK_D_T dut(S, R, clk, rst, Q_jk, Q_d, Q_t);
initial begin 
        clk = 0;
       forever #5 clk = ~clk;
       end 
       
 initial begin
        rst=1;
        S = 0;
        R = 0;
        #10;
        rst=0;
    end
    
    always begin
        S=0;
        R=0;
        #10;
        S=0;
        R=1;
        #10;
        S=1;
        R=0;
        #10;
        S=1;
        R=1;
        #10;

    end
  initial begin
  $dumpfile("test_bench.vcd");
  $dumpvars(0,test_bench);
  $monitor("\t clk: %d  S: %d  R: %d  Q_jk: %d  Q_d: %d  Q_t:%d", clk,S,R,Q_jk, Q_d, Q_t);
  #90 $finish;
  end
endmodule


module D_flipflop(
input clk,reset,d,
output reg Q);

always@(posedge clk) begin 
if({reset}) Q<=1'b0;
else 
Q<=d; 

end
endmodule 